module example(input x, output y);
   

always_ff @(posedge clk)
begin
   a <= b;
end

